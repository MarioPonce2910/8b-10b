module serialization(clk,rst,data_in,data_out);
    input clk,rst;
    input [7:0] data_in;
    output [9:0] data_out;
    wire flag;
        reg [5:0] 5b/6b [31:0] [1:0];
        reg [3:0] 3b/4b [7:0] [1:0];

            initial begin
            //0
                5b/6b [0] [0] = 6'b100111; 
                5b/6b [0] [1] = 6'b011000;
            //1
                5b/6b [1] [0] = 6'b011101; 
                5b/6b [1] [1] = 6'b100010;
            //2
                5b/6b [2] [0] = 6'b101101; 
                5b/6b [2] [1] = 6'b010010;
            //3
                5b/6b [3] [0] = 6'b110001; 
                5b/6b [3] [1] = 6'b110001;
            //4
                5b/6b [4] [0] = 6'b110101; 
                5b/6b [4] [1] = 6'b001010;
            //5
                5b/6b [5] [0] = 6'b101001; 
                5b/6b [5] [1] = 6'b101001;
            //6
                5b/6b [6] [0] = 6'b011001; 
                5b/6b [6] [1] = 6'b011001;
            //7
                5b/6b [7] [0] = 6'b111000; 
                5b/6b [7] [1] = 6'b000111;
            //8
                5b/6b [8] [0] = 6'b111001; 
                5b/6b [8] [1] = 6'b000101;
            //9
                5b/6b [9] [0] = 6'b100101; 
                5b/6b [9] [1] = 6'b100101;
            //10
                5b/6b [10] [0] = 6'b010101; 
                5b/6b [10] [1] = 6'b010101;
            //11
                5b/6b [11] [0] = 6'b110100; 
                5b/6b [11] [1] = 6'b110100;
            //12
                5b/6b [12] [0] = 6'b001101; 
                5b/6b [12] [1] = 6'b001101;
            //13
                5b/6b [13] [0] = 6'b101100; 
                5b/6b [13] [1] = 6'b101100;
            //14
                5b/6b [14] [0] = 6'b011100; 
                5b/6b [14] [1] = 6'b011100;
            //15
                5b/6b [15] [0] = 6'b010111; 
                5b/6b [15] [1] = 6'b101000;
            //16
                5b/6b [16] [0] = 6'b011011; 
                5b/6b [16] [1] = 6'b100100;
            //17
                5b/6b [17] [0] = 6'b100011; 
                5b/6b [17] [1] = 6'b100011;
            //18
                5b/6b [18] [0] = 6'b010011; 
                5b/6b [18] [1] = 6'b010011;
            //19
                5b/6b [19] [0] = 6'b110010; 
                5b/6b [19] [1] = 6'b110010;
            //20
                5b/6b [20] [0] = 6'b001011; 
                5b/6b [20] [1] = 6'b001011;
            //21
                5b/6b [21] [0] = 6'b101010; 
                5b/6b [21] [1] = 6'b101010;
            //22
                5b/6b [22] [0] = 6'b011010; 
                5b/6b [22] [1] = 6'b011010;
            //23
                5b/6b [23] [0] = 6'b111010; 
                5b/6b [23] [1] = 6'b000101;
            //24
                5b/6b [24] [0] = 6'b110011; 
                5b/6b [24] [1] = 6'b001100;
            //25
                5b/6b [25] [0] = 6'b100110; 
                5b/6b [25] [1] = 6'b100110;
            //26
                5b/6b [26] [0] = 6'b010110; 
                5b/6b [26] [1] = 6'b010110;
            //27
                5b/6b [27] [0] = 6'b110110; 
                5b/6b [27] [1] = 6'b001001;
            //28
                5b/6b [28] [0] = 6'b001110; 
                5b/6b [28] [1] = 6'b001110;
            //29
                5b/6b [29] [0] = 6'b101110; 
                5b/6b [29] [1] = 6'b010001;
            //30
                5b/6b [30] [0] = 6'b011110; 
                5b/6b [30] [1] = 6'b100001;
            //31
                5b/6b [31] [0] = 6'b; 
                5b/6b [31] [1] = 6'b100010;
            end

    always@(posedge clk)
        begin
            if(flag == 1)
                begin
                    for ( = ; ; ) begin
                        
                    end
                end
        end




endmodule